module hello_world_in_verilog;
initial 
  begin
    $display ("Hello World");
    $finish;
  end
endmodule